// jeden modul RAM z paramterami.

module ram#(
    parameter
)
(
    input wire clk
);



endmodule