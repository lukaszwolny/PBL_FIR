////////////////////////////////////////////////////////////////////////
//   główny moduł dla AXI.
//   Do testów w cocoTB
///////////////////////////////////////////////////////////////////////

//AXI

//MUX'y
//MUX_AXI_wej

//MUX_AXI_wyj

//RAM (wej)

//RAM (wyj)
